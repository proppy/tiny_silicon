module tiny_user_project (vccd1,
    vssd1,
    io_in,
    io_oeb,
    io_out);
 input vccd1;
 input vssd1;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire net48;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net49;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net50;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net18;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net19;
 wire net38;
 wire net39;
 wire net20;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire \mod.flipflop1.clk ;
 wire \mod.flipflop1.d ;
 wire \mod.flipflop3.d ;
 wire \mod.flipflop4.d ;
 wire \mod.flipflop5.d ;
 wire \mod.flipflop6.d ;
 wire \mod.flop2.clk ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;

 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _009_ (.A1(net3),
    .A2(net2),
    .B(net1),
    .ZN(_000_),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _010_ (.I(_000_),
    .ZN(\mod.flop2.clk ),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _011_ (.I(net2),
    .ZN(_001_),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _012_ (.I(_001_),
    .Z(_002_),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _013_ (.I(net1),
    .ZN(_003_),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _014_ (.A1(net3),
    .A2(_002_),
    .B(_003_),
    .ZN(\mod.flipflop1.clk ),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _015_ (.A1(_002_),
    .A2(net5),
    .Z(_004_),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _016_ (.I(_004_),
    .Z(\mod.flipflop3.d ),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _017_ (.A1(_002_),
    .A2(net4),
    .Z(_005_),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _018_ (.I(_005_),
    .Z(\mod.flipflop1.d ),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _019_ (.A1(_002_),
    .A2(net8),
    .Z(_006_),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _020_ (.I(_006_),
    .Z(\mod.flipflop6.d ),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _021_ (.A1(_001_),
    .A2(net7),
    .Z(_007_),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _022_ (.I(_007_),
    .Z(\mod.flipflop5.d ),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _023_ (.A1(_001_),
    .A2(net6),
    .Z(_008_),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _024_ (.I(_008_),
    .Z(\mod.flipflop4.d ),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _025_ (.D(\mod.flipflop1.d ),
    .CLK(\mod.flipflop1.clk ),
    .Q(net9),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _026_ (.D(\mod.flipflop1.d ),
    .CLK(\mod.flop2.clk ),
    .Q(net14),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _027_ (.D(\mod.flipflop3.d ),
    .CLK(\mod.flipflop1.clk ),
    .Q(net10),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _028_ (.D(\mod.flipflop3.d ),
    .CLK(\mod.flop2.clk ),
    .Q(net15),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _029_ (.D(\mod.flipflop4.d ),
    .CLK(\mod.flipflop1.clk ),
    .Q(net11),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _030_ (.D(\mod.flipflop4.d ),
    .CLK(\mod.flop2.clk ),
    .Q(net16),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _031_ (.D(\mod.flipflop5.d ),
    .CLK(\mod.flipflop1.clk ),
    .Q(net12),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _032_ (.D(\mod.flipflop6.d ),
    .CLK(\mod.flipflop1.clk ),
    .Q(net13),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_18 (.ZN(net18),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_19 (.ZN(net19),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_20 (.ZN(net20),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_21 (.ZN(net21),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_22 (.ZN(net22),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_23 (.ZN(net23),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_24 (.ZN(net24),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_25 (.ZN(net25),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_26 (.ZN(net26),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_27 (.ZN(net27),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_28 (.ZN(net28),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_29 (.ZN(net29),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_30 (.ZN(net30),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_31 (.ZN(net31),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_32 (.ZN(net32),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_33 (.ZN(net33),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_34 (.ZN(net34),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_35 (.ZN(net35),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_36 (.ZN(net36),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_37 (.ZN(net37),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_38 (.ZN(net38),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_39 (.ZN(net39),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_40 (.ZN(net40),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_41 (.ZN(net41),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_42 (.ZN(net42),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_43 (.ZN(net43),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_44 (.ZN(net44),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_45 (.ZN(net45),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_46 (.ZN(net46),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_47 (.ZN(net47),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_48 (.ZN(net48),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_49 (.ZN(net49),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_50 (.ZN(net50),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_51 (.ZN(net51),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_52 (.ZN(net52),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_53 (.ZN(net53),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_54 (.ZN(net54),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_55 (.ZN(net55),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_56 (.ZN(net56),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_57 (.ZN(net57),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_58 (.ZN(net58),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_59 (.ZN(net59),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_60 (.ZN(net60),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_61 (.ZN(net61),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_62 (.ZN(net62),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_63 (.ZN(net63),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_64 (.ZN(net64),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_65 (.ZN(net65),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_66 (.ZN(net66),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_67 (.ZN(net67),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_68 (.ZN(net68),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_69 (.ZN(net69),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_70 (.ZN(net70),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_71 (.ZN(net71),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_72 (.ZN(net72),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_73 (.ZN(net73),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_74 (.ZN(net74),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_75 (.ZN(net75),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_76 (.ZN(net76),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_77 (.ZN(net77),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_78 (.ZN(net78),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_79 (.ZN(net79),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_80 (.ZN(net80),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_81 (.ZN(net81),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_82 (.ZN(net82),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_83 (.ZN(net83),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_84 (.ZN(net84),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__019__A1 (.I(_002_),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_110 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_111 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_112 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_113 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_114 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_115 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_116 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_117 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_118 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_119 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_120 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_121 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_122 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_123 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_124 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_125 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_126 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_127 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_128 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_129 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_130 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_131 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_132 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_133 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_134 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_135 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_136 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_138 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_139 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_140 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_142 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_143 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_145 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_146 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_147 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_148 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_149 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_150 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_151 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_152 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_153 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_154 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_155 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_156 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_157 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_158 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_159 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_160 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_161 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_162 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_163 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_164 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_165 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_166 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_167 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_168 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_169 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_170 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_171 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_173 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_174 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_175 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_177 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_178 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_180 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_181 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_182 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_183 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_184 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_185 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_186 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_187 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_188 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_189 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_190 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_191 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_192 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_193 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_194 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_195 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_196 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_197 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_198 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_199 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_200 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_201 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_202 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_203 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_204 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_205 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_206 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_207 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_209 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_210 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_211 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_288 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_289 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(io_in[12]),
    .Z(net1),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(io_in[13]),
    .Z(net2),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(io_in[14]),
    .Z(net3),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(io_in[15]),
    .Z(net4),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(io_in[16]),
    .Z(net5),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(io_in[17]),
    .Z(net6),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(io_in[18]),
    .Z(net7),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(io_in[19]),
    .Z(net8),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output9 (.I(net9),
    .Z(io_out[20]),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output10 (.I(net10),
    .Z(io_out[21]),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output11 (.I(net11),
    .Z(io_out[22]),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output12 (.I(net12),
    .Z(io_out[23]),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output13 (.I(net13),
    .Z(io_out[24]),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output14 (.I(net14),
    .Z(io_out[25]),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output15 (.I(net15),
    .Z(io_out[26]),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output16 (.I(net16),
    .Z(io_out[27]),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_17 (.ZN(net17),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__017__A1 (.I(_002_),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__015__A1 (.I(_002_),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__014__A2 (.I(_002_),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[12]),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[13]),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[14]),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[15]),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[16]),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[17]),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[18]),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[19]),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__011__I (.I(net2),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__009__A2 (.I(net2),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__014__A1 (.I(net3),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__009__A1 (.I(net3),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__017__A2 (.I(net4),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__015__A2 (.I(net5),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__023__A2 (.I(net6),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__021__A2 (.I(net7),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__019__A2 (.I(net8),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output9_I (.I(net9),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output11_I (.I(net11),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output12_I (.I(net12),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output13_I (.I(net13),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output14_I (.I(net14),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output15_I (.I(net15),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output16_I (.I(net16),
    .VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_190 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_192 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_197 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_205 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_220 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_222 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_227 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_252 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_268 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_270 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_275 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_282 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_298 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_300 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_305 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_309 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_311 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_325 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_335 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_343 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_347 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_352 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_365 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_371 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_383 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_387 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_395 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_401 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_411 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_7 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_13 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_45 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_61 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_69 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_409 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_416 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_412 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_414 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_7 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_412 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_414 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_7 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_412 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_414 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_7 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_416 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_412 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_414 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_7 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_23 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_31 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_416 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_7 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_23 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_31 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_416 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_7 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_23 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_31 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_412 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_414 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_7 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_23 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_31 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_416 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_416 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_7 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_412 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_414 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_17 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_21 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_53 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_69 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_412 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_414 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_7 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_416 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_7 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_23 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_31 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_412 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_414 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_7 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_23 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_31 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_416 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_7 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_23 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_31 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_416 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_412 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_414 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_7 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_23 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_31 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_416 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_412 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_414 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_7 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_412 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_414 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_7 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_412 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_414 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_7 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_140 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_156 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_158 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_163 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_167 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_171 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_175 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_416 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_148 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_150 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_159 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_161 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_170 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_174 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_178 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_210 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_124 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_128 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_132 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_142 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_173 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_416 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_121 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_129 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_133 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_174 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_182 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_190 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_206 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_210 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_7 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_23 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_31 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_116 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_120 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_123 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_131 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_172 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_188 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_196 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_200 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_232 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_416 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_5 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_69 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_121 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_131 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_147 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_162 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_193 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_209 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_350 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_411 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_17 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_21 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_29 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_33 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_108 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_124 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_132 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_136 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_139 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_145 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_179 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_209 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_241 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_245 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_250 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_321 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_385 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_392 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_408 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_416 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_7 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_13 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_19 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_51 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_67 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_144 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_148 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_153 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_161 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_192 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_208 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_215 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_286 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_294 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_300 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_332 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_348 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_352 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_357 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_389 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_405 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_413 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_417 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_419 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_9 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_15 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_19 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_37 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_40 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_48 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_52 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_54 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_59 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_67 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_69 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_72 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_77 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_85 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_89 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_97 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_107 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_112 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_128 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_132 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_134 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_139 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_142 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_173 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_177 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_192 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_198 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_206 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_212 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_228 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_233 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_241 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_247 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_255 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_259 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_263 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_271 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_275 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_279 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_282 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_297 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_299 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_314 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_317 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_329 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_337 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_341 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_347 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_349 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_352 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_360 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_364 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_368 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_384 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_387 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_403 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_411 (.VDD(vccd1),
    .VSS(vssd1));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_419 (.VDD(vccd1),
    .VSS(vssd1));
 assign io_oeb[0] = net47;
 assign io_oeb[10] = net57;
 assign io_oeb[11] = net58;
 assign io_oeb[12] = net59;
 assign io_oeb[13] = net60;
 assign io_oeb[14] = net61;
 assign io_oeb[15] = net62;
 assign io_oeb[16] = net63;
 assign io_oeb[17] = net64;
 assign io_oeb[18] = net65;
 assign io_oeb[19] = net66;
 assign io_oeb[1] = net48;
 assign io_oeb[20] = net67;
 assign io_oeb[21] = net68;
 assign io_oeb[22] = net69;
 assign io_oeb[23] = net70;
 assign io_oeb[24] = net71;
 assign io_oeb[25] = net72;
 assign io_oeb[26] = net73;
 assign io_oeb[27] = net74;
 assign io_oeb[28] = net75;
 assign io_oeb[29] = net76;
 assign io_oeb[2] = net49;
 assign io_oeb[30] = net77;
 assign io_oeb[31] = net78;
 assign io_oeb[32] = net79;
 assign io_oeb[33] = net80;
 assign io_oeb[34] = net81;
 assign io_oeb[35] = net82;
 assign io_oeb[36] = net83;
 assign io_oeb[37] = net84;
 assign io_oeb[3] = net50;
 assign io_oeb[4] = net51;
 assign io_oeb[5] = net52;
 assign io_oeb[6] = net53;
 assign io_oeb[7] = net54;
 assign io_oeb[8] = net55;
 assign io_oeb[9] = net56;
 assign io_out[0] = net17;
 assign io_out[10] = net27;
 assign io_out[11] = net28;
 assign io_out[12] = net29;
 assign io_out[13] = net30;
 assign io_out[14] = net31;
 assign io_out[15] = net32;
 assign io_out[16] = net33;
 assign io_out[17] = net34;
 assign io_out[18] = net35;
 assign io_out[19] = net36;
 assign io_out[1] = net18;
 assign io_out[28] = net37;
 assign io_out[29] = net38;
 assign io_out[2] = net19;
 assign io_out[30] = net39;
 assign io_out[31] = net40;
 assign io_out[32] = net41;
 assign io_out[33] = net42;
 assign io_out[34] = net43;
 assign io_out[35] = net44;
 assign io_out[36] = net45;
 assign io_out[37] = net46;
 assign io_out[3] = net20;
 assign io_out[4] = net21;
 assign io_out[5] = net22;
 assign io_out[6] = net23;
 assign io_out[7] = net24;
 assign io_out[8] = net25;
 assign io_out[9] = net26;
endmodule
